-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Sat Sep 28 21:59:47 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY \7_seg_driver\ IS 
	PORT
	(
		D0 :  IN  STD_LOGIC;
		D1 :  IN  STD_LOGIC;
		D2 :  IN  STD_LOGIC;
		D3 :  IN  STD_LOGIC;
		Ripple_Blanking :  IN  STD_LOGIC;
		Seg_0 :  OUT  STD_LOGIC;
		Seg_1 :  OUT  STD_LOGIC;
		Seg_2 :  OUT  STD_LOGIC;
		Seg_3 :  OUT  STD_LOGIC;
		Seg_4 :  OUT  STD_LOGIC;
		Seg_5 :  OUT  STD_LOGIC;
		Seg_6 :  OUT  STD_LOGIC;
		Ripple_Blanking_Carry :  OUT  STD_LOGIC
	);
END \7_seg_driver\;

ARCHITECTURE bdf_type OF \7_seg_driver\ IS 

SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;


BEGIN 
Ripple_Blanking_Carry <= SYNTHESIZED_WIRE_89;



SYNTHESIZED_WIRE_67 <= SYNTHESIZED_WIRE_86 AND SYNTHESIZED_WIRE_87 AND SYNTHESIZED_WIRE_88 AND D0;


SYNTHESIZED_WIRE_11 <= D3 OR D1 OR D0 OR D2;


Seg_0 <= SYNTHESIZED_WIRE_89 OR SYNTHESIZED_WIRE_4;


Seg_1 <= SYNTHESIZED_WIRE_89 OR SYNTHESIZED_WIRE_6;


Seg_2 <= SYNTHESIZED_WIRE_89 OR SYNTHESIZED_WIRE_8;


Seg_3 <= SYNTHESIZED_WIRE_89 OR SYNTHESIZED_WIRE_10;


SYNTHESIZED_WIRE_21 <= NOT(SYNTHESIZED_WIRE_11);



Seg_4 <= SYNTHESIZED_WIRE_89 OR SYNTHESIZED_WIRE_13;


Seg_5 <= SYNTHESIZED_WIRE_89 OR SYNTHESIZED_WIRE_15;


Seg_6 <= SYNTHESIZED_WIRE_89 OR SYNTHESIZED_WIRE_17;


SYNTHESIZED_WIRE_66 <= SYNTHESIZED_WIRE_86 AND D2 AND SYNTHESIZED_WIRE_88 AND SYNTHESIZED_WIRE_90;


SYNTHESIZED_WIRE_89 <= SYNTHESIZED_WIRE_21 AND Ripple_Blanking;


SYNTHESIZED_WIRE_69 <= SYNTHESIZED_WIRE_86 AND D2 AND SYNTHESIZED_WIRE_88 AND D0;


SYNTHESIZED_WIRE_68 <= SYNTHESIZED_WIRE_86 AND D2 AND D1 AND SYNTHESIZED_WIRE_90;


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_86 AND SYNTHESIZED_WIRE_87 AND D1 AND SYNTHESIZED_WIRE_90;


SYNTHESIZED_WIRE_79 <= SYNTHESIZED_WIRE_86 AND SYNTHESIZED_WIRE_87 AND SYNTHESIZED_WIRE_88 AND D0;


SYNTHESIZED_WIRE_77 <= SYNTHESIZED_WIRE_86 AND D2 AND SYNTHESIZED_WIRE_88 AND SYNTHESIZED_WIRE_90;


SYNTHESIZED_WIRE_78 <= SYNTHESIZED_WIRE_86 AND D2 AND D1 AND D0;


SYNTHESIZED_WIRE_80 <= D3 AND SYNTHESIZED_WIRE_87 AND SYNTHESIZED_WIRE_88 AND D0;


SYNTHESIZED_WIRE_82 <= SYNTHESIZED_WIRE_86 AND SYNTHESIZED_WIRE_87 AND SYNTHESIZED_WIRE_88 AND D0;


SYNTHESIZED_WIRE_81 <= SYNTHESIZED_WIRE_86 AND SYNTHESIZED_WIRE_87 AND D1 AND D0;


SYNTHESIZED_WIRE_86 <= NOT(D3);



SYNTHESIZED_WIRE_83 <= SYNTHESIZED_WIRE_86 AND D2 AND SYNTHESIZED_WIRE_88 AND D0;


SYNTHESIZED_WIRE_84 <= SYNTHESIZED_WIRE_86 AND D2 AND D1 AND D0;


SYNTHESIZED_WIRE_85 <= SYNTHESIZED_WIRE_86 AND D2 AND SYNTHESIZED_WIRE_88 AND SYNTHESIZED_WIRE_90;


SYNTHESIZED_WIRE_70 <= SYNTHESIZED_WIRE_86 AND SYNTHESIZED_WIRE_87 AND SYNTHESIZED_WIRE_88 AND D0;


SYNTHESIZED_WIRE_73 <= SYNTHESIZED_WIRE_86 AND SYNTHESIZED_WIRE_87 AND D1 AND SYNTHESIZED_WIRE_90;


SYNTHESIZED_WIRE_71 <= SYNTHESIZED_WIRE_86 AND SYNTHESIZED_WIRE_87 AND D1 AND D0;


SYNTHESIZED_WIRE_72 <= SYNTHESIZED_WIRE_86 AND D2 AND D1 AND D0;


SYNTHESIZED_WIRE_76 <= SYNTHESIZED_WIRE_86 AND SYNTHESIZED_WIRE_87 AND SYNTHESIZED_WIRE_88 AND SYNTHESIZED_WIRE_90;


SYNTHESIZED_WIRE_74 <= SYNTHESIZED_WIRE_86 AND SYNTHESIZED_WIRE_87 AND SYNTHESIZED_WIRE_88 AND D0;


SYNTHESIZED_WIRE_75 <= SYNTHESIZED_WIRE_86 AND D0 AND D1 AND D2;


SYNTHESIZED_WIRE_87 <= NOT(D2);



SYNTHESIZED_WIRE_4 <= SYNTHESIZED_WIRE_66 OR SYNTHESIZED_WIRE_67;


SYNTHESIZED_WIRE_6 <= SYNTHESIZED_WIRE_68 OR SYNTHESIZED_WIRE_69;


SYNTHESIZED_WIRE_15 <= SYNTHESIZED_WIRE_70 OR SYNTHESIZED_WIRE_71 OR SYNTHESIZED_WIRE_72 OR SYNTHESIZED_WIRE_73;


SYNTHESIZED_WIRE_17 <= SYNTHESIZED_WIRE_74 OR SYNTHESIZED_WIRE_75 OR SYNTHESIZED_WIRE_76;


SYNTHESIZED_WIRE_10 <= SYNTHESIZED_WIRE_77 OR SYNTHESIZED_WIRE_78 OR SYNTHESIZED_WIRE_79;


SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_80 OR SYNTHESIZED_WIRE_81 OR SYNTHESIZED_WIRE_82 OR SYNTHESIZED_WIRE_83 OR SYNTHESIZED_WIRE_84 OR SYNTHESIZED_WIRE_85;


SYNTHESIZED_WIRE_88 <= NOT(D1);



SYNTHESIZED_WIRE_90 <= NOT(D0);



END bdf_type;